module testbench();
    reg in;
    wire out;
    not test_unit(in,out);

    initial begin

    end
endmodule