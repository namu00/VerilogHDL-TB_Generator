module t_latch(t, out);
    input t;
    output out;

    /* */

endmodule