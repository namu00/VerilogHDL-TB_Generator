module d_latch(d, out);
    input d;
    output out;

    assign out = d;
endmodule